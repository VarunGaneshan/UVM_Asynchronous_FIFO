`define ADDR_WIDTH 4
`define DATA_WIDTH 8
`define WCLK_PERIOD 10
`define RCLK_PERIOD 20
`define FIFO_DEPTH (1<<`ADDR_WIDTH)

`define NUM_WRITE_TRANS_WR `FIFO_DEPTH+6+9
`define NUM_READ_TRANS_WR `FIFO_DEPTH+6+8

`define NUM_WRITE_TRANS_WTR `FIFO_DEPTH+2
`define NUM_READ_LOW_WTR (`FIFO_DEPTH/2)+1
`define NUM_READ_TRANS_WTR `FIFO_DEPTH+1