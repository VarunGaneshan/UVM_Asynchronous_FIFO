`define ADDR_WIDTH 4
`define DATA_WIDTH 8
`define WCLK_PERIOD 10
`define RCLK_PERIOD 20
`define FIFO_DEPTH (1<<`ADDR_WIDTH)
`define NUM_WRITE_TRANS `FIFO_DEPTH+6+10
`define NUM_READ_TRANS `FIFO_DEPTH+6+9